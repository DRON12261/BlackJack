.   3   f&  5   e&  A   `&  Q   f&  4   c&  K   `&  X   e&  2   c&  8   `&  8   f&  Q   c&  6   e&  K   f&  9   c&  6   `&  6   f&  7   f&  J   c&  7   e&  J   `&  K   e&  J   e&  5   c&  5   f&  3   c&  8   e&  A   f&  9   f&  9   e&  3   `&  Q   e&  8   c&  6   c&  7   `&  A   e&  4   e&  K   c&  4   `&  4   f&  5   `&  X   `&  9   `&  Q   `&  A   c&  2   f&  X   f&     12312       2   e&  X   c&            1243      3   e&  J   f&                    
Дилер   2   `&  7   c&                       